// Code your design here
module or_gate(y,a,b);
input a,b;
output reg y;
assign y=a|b;
endmodule;