// Code your design here
module and_gate(a,b,y);
input a,b;
output reg y;
assign y=a&b;
endmodule;
